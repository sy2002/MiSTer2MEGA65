// Taken from MiSTer's sys/sys_top.v @ 390f45a by sy2002 in May 2023
//
// CSync generation
// Shifts HSync left by 1 HSync period during VSync

module csync
(
    input  clk,
    input  hsync,
    input  vsync,

    output csync
);

assign csync = (csync_vs ^ csync_hs);

reg csync_hs, csync_vs;
always @(posedge clk) begin
    reg prev_hs;
    reg [15:0] h_cnt, line_len, hs_len;

    // Count line/Hsync length
    h_cnt <= h_cnt + 1'd1;

    prev_hs <= hsync;
    if (prev_hs ^ hsync) begin
        h_cnt <= 0;
        if (hsync) begin
            line_len <= h_cnt - hs_len;
            csync_hs <= 0;
        end
        else hs_len <= h_cnt;
    end
    
    if (~vsync) csync_hs <= hsync;
    else if(h_cnt == line_len) csync_hs <= 1;
    
    csync_vs <= vsync;
end

endmodule
